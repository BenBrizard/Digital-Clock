-------------------------------------------------------------------------------
-- Title      : ROM_data
-- Project    : Horloge numerique - projet 3 ELE3311 - hiver 2019
-------------------------------------------------------------------------------
-- File       : ROM_data.vhd
-- Author     : AR
-- Created    : 2019-03-03
-- Last update: 2019-03-09
-------------------------------------------------------------------------------
-- Description: ROM contenant les commandes et les caractères à dessiner sur
--              l'écran OLED. 
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package ROM_data is

type ROM_cmd_t is array (0 to 511) of std_logic_vector(63 downto 0);
constant CMD_MEM : ROM_cmd_t := (
--X"ffffff0100138800", X"ffffff40000000AE", X"ffffff1000138800", X"ffffff3000138800", X"ffffff400000008D", X"ffffff4000000014", X"ffffff40000000D9", X"ffffff40000000F1",         --power on sequence
--X"ffffff0407A12000", X"ffffff4000000081", X"ffffff400000000F", X"ffffff40000000A0", X"ffffff40000000C0", X"ffffff40000000DA", X"ffffff4000000000", X"ffffff40000000AF",
X"ffffff0100000200", X"ffffff40000000AE", X"ffffff1000000200", X"ffffff3000000200", X"ffffff400000008D", X"ffffff4000000014", X"ffffff40000000D9", X"ffffff40000000F1",       --simulation power on
X"ffffff0400000200", X"ffffff4000000081", X"ffffff400000000F", X"ffffff40000000A0", X"ffffff40000000C0", X"ffffff40000000DA", X"ffffff4000000000", X"ffffffC0000000AF",
X"ffffff4000000020", X"ffffffC000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff40000000AE", X"ffffff0C07A12000", X"ffffff8300138800", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",         --power off sequence           
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000",
X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000", X"ffffff0000000000"
);

type ROM_char_t is array (0 to 1023) of std_logic_vector(7 downto 0);
constant CHAR_MEM : ROM_char_t := (
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","11111100","11111100","00000011","00000011","00000011","00000011","00000011","00000011","11111100","11111100","00000000","00000000","00000000",
"00000000","00000000","00000000","00111111","00111111","11000000","11000000","11000000","11000000","11000000","11000000","00111111","00111111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00001100","00001100","11111111","11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","11000000","11000000","11111111","11111111","11000000","11000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00001100","00001100","00000011","00000011","00000011","00000011","11000011","11000011","00111100","00111100","00000000","00000000","00000000",
"00000000","00000000","00000000","11110000","11110000","11001100","11001100","11000011","11000011","11000000","11000000","11000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00001100","00001100","00000011","00000011","11000011","11000011","11000011","11000011","00111100","00111100","00000000","00000000","00000000",
"00000000","00000000","00000000","01100000","01100000","11000000","11000000","11000000","11000000","11000000","11000000","00111111","00111111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","11000000","11000000","00110000","00110000","00001100","00001100","11111111","11111111","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000011","00000011","00000011","00000011","00000011","00000011","11111111","11111111","00000011","00000011","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","11111111","11111111","11000011","11000011","11000011","11000011","11000011","00000011","00000011","00000000","00000000","00000000",
"00000000","00000000","00000000","00110000","00110000","11000000","11000000","11000000","11000000","11000000","11000000","00111111","00111111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","11110000","11110000","11001100","11001100","11000011","11000011","11000011","11000011","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00111111","00111111","11000000","11000000","11000000","11000000","11000000","11000000","00111111","00111111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000011","00000011","00000011","00000011","00000011","00000011","11110011","11110011","00001111","00001111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","11110000","11110000","00001111","00001111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00111100","00111100","11000011","11000011","11000011","11000011","11000011","11000011","00111100","00111100","00000000","00000000","00000000",
"00000000","00000000","00000000","00111111","00111111","11000000","11000000","11000000","11000000","11000000","11000000","00111111","00111111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","11111100","11111100","00000011","00000011","00000011","00000011","00000011","00000011","11111100","11111100","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","11000011","11000011","11000011","11000011","00110011","00110011","00001111","00001111","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00111100","00111100","00111100","00111100","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00111100","00111100","00111100","00111100","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","11111111","11111111","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
"00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000"
);

end package ROM_data;
